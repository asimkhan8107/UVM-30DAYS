
`include "interface.sv"
`include "sequence_item.sv"
`include "dff.v"
`include "sequences.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor_in.sv"
`include "agent1.sv"
`include "monitor_out.sv"
`include "agent2.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"